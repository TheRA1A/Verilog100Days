module test1 ();

endmodule
